package shared_pkg;
	
	bit test_finished;

	int c_count_ALURes, c_count_PCNext, c_count_RD_m, c_count_MemWr, c_count_MemRd, c_count_Stall;
    int e_count_ALURes, e_count_PCNext, e_count_RD_m, e_count_MemWr, e_count_MemRd, e_count_Stall;

endpackage